`define RISCV_FORMAL
`define RISCV_FORMAL_NRET 1
`define RISCV_FORMAL_XLEN 32
`define RISCV_FORMAL_ILEN 32
`define RISCV_FORMAL_CHECKER rvfi_reg_check
`define RISCV_FORMAL_RESET_CYCLES 15
`define RISCV_FORMAL_CHECK_CYCLE 25
`define RISCV_FORMAL_CHANNEL_IDX 0
`define RISCV_FORMAL_ALIGNED_MEM
`define RISCV_FORMAL_ALTOPS
`include "rvfi_macros.vh"
